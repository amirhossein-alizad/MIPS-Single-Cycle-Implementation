`timescale 1ns/1ns
module adder(input [31:0] inp1, inp2, output  [31:0]  out);
  assign out = inp1 + inp2;
endmodule

